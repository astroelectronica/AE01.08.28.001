.title KiCad schematic
.include "models/LUXEON_Rebel_ES_H_and_5630_diode_models.txt"
D3 /IN /1 LXML-PWN2-VFBin_R
V1 /IN 0 {VIN}
D4 /IN /1 LXML-PWN2-VFBin_R
D1 /IN /1 LXML-PWN2-VFBin_R
D2 /IN /1 LXML-PWN2-VFBin_R
D7 /1 /2 LXML-PWN2-VFBin_R
D8 /1 /2 LXML-PWN2-VFBin_R
D5 /1 /2 LXML-PWN2-VFBin_R
D6 /1 /2 LXML-PWN2-VFBin_R
D11 /2 /3 LXML-PWN2-VFBin_R
D12 /2 /3 LXML-PWN2-VFBin_R
D9 /2 /3 LXML-PWN2-VFBin_R
D10 /2 /3 LXML-PWN2-VFBin_R
D15 /3 0 LXML-PWN2-VFBin_R
D16 /3 0 LXML-PWN2-VFBin_R
D13 /3 0 LXML-PWN2-VFBin_R
D14 /3 0 LXML-PWN2-VFBin_R
.end
